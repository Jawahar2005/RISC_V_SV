`include "packet.sv"
`include "interface.sv"
`include "clock_generation.sv"
`include "alu_random_test.sv"
`include "alu_unit_test.sv"
`include "alu_edgecase_test.sv"
`include "instruction_memory_test.sv"
`include "reg_file_random_test.sv"
`include "reg_file_read_test.sv"
`include "reg_file_write_test.sv"
`include "reg_file_disable_write_test.sv"
`include "control_unit_test.sv"
`include "control_unit_random_test.sv"
`include "alu_control_unit_test.sv"
`include "data_memory_test.sv"
`include "data_memory_write_test.sv"
`include "data_memory_read_test.sv"
`include "data_memory_disable_read_test.sv"
`include "data_memory_disable_write_test.sv"
