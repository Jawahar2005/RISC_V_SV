`ifndef PARAMETER_H_
`define PARAMETER_H_
`define col 16 
`define row_i 15 
`define row_d 8  
`define filename "test.data"
`define simulation_time #160
`endif
